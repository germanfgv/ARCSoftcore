
// SharkBoad SystemModule
//
// Top Level Design for the Xilinx Spartan 3-100E Device
//---------------------------------------------------------------------------

/*#
# SharkBoad
# Copyright (C) 2012 Bogotá, Colombia
#
# This program is free software: you can redistribute it and/or modify
# it under the terms of the GNU General Public License as published by
# the Free Software Foundation, version 3 of the License.
#
# This program is distributed in the hope that it will be useful,
# but WITHOUT ANY WARRANTY; without even the implied warranty of
# MERCHANTABILITY or FITNESS FOR A PARTICULAR PURPOSE.  See the
# GNU General Public License for more details.
#
# You should have received a copy of the GNU General Public License
# along with this program.  If not, see <http://www.gnu.org/licenses/>.
#*/

module system
#(parameter	clk_freq	= 50000000) 
(
	input		clk, rst, rx,
	output		tx,useless,full


);
/*Declaración de cables*/

	wire [7:0] w_edata;	

/*Decaración demódulos*/

	/*Control section: Esté módulo cnntrola la operación del datapath. 
	Contiene toda la lógica que permite decidir 
        los pasos a seguir para llevar a cabo la intrucciónes de la Main Memory.*/

	uart uart_echo(
	    	.clk(clk), 
		.reset(rst),
	    	.rd_uart(~w_empty),
		.wr_uart(~w_empty), 
		.rx(rx),
	    	.w_data(w_edata), 
	    	.tx_full(full), 
		.rx_empty(w_empty), 
		.tx(tx),
	    	.r_data(w_edata),
	    	.useless(useless)
	);




endmodule
