module reset(
/*Este ódulo se encarga de devolver la MIR (y en general toda la control section) a un estado inicial en el momento en que una señal de rst entra al sistema*/
);

