module control_store (
input rst,
input [10:0]	address,
output reg[40:0] mir 
);




always@(*)
begin

if (rst)
	mir=41'b10000001000000100101010010100000000000000;	
else
begin
	case(address)
0:mir=41'b10000001000000100101010010100000000000000;//Initial instruction
1:mir=41'b00000000000000000000000010111100000000000;//DECODE
1152:mir=41'b10010100000000000000100101011011111111111;//sethi (Lshift of ri to a chossen register)

/*call*/
1280:mir=41'b10000001000000001111000010100000000000000;//pc to R15
1281:mir=41'b10010101001010100001000100000000000000000;//left-shift of ri  to temp0
1282:mir=41'b10000101000010100001000100000000000000000;// left-shift of temp0 to temp0
1283:mir=41'b10000001000010100000000100011000000000000;// new pc: adding pc and temp0
1600:mir=41'b00000000000000000000000010110111001000010;
1601:mir=41'b00000010000001000000100001111011111111111;
1602:mir=41'b10010100000000100001000110000000000000000;
1603:mir=41'b00000011000010000000100001111011111111111;
1604:mir=41'b00000000000000000000000010110111001000110;
1605:mir=41'b00000010000001000000100000011011111111111;
1606:mir=41'b10010100000000100001000101100000000000000;
1607:mir=41'b00000011000010000000100000011011111111111;
1608:mir=41'b00000000000000000000000010110111001001010;
1609:mir=41'b00000010000001000000100000111011111111111;
1610:mir=41'b10010100000000100001000101100000000000000;
1611:mir=41'b00000011000010000000100000111011111111111;
1624:mir=41'b00000000000000000000000010110111001011010;
1625:mir=41'b00000010000001000000100001011011111111111;
1626:mir=41'b10010100000000100001000101100000000000000;
1627:mir=41'b00000011000010000000100001011011111111111;
1688:mir=41'b00000000000000000000000010100011010011010;
1689:mir=41'b00000010000001000000100010011011111111111;
1690:mir=41'b10010100000000100001000101100000000000000;
1691:mir=41'b00000011000010000000100010011011111111111;
1760:mir=41'b00000000000000000000000010110111011100010;
1761:mir=41'b00000010000001100000000100011000000000000;
1762:mir=41'b10010100000000100001000110000000000000000;
1763:mir=41'b00000011000010100000000100011000000000000;
1792:mir=41'b00000010000001100001000100010111100000010;

1793:mir=41'b10000101000010000000110010111011111111111;
1794:mir=41'b10010100000000100001000110000000000000000;
1795:mir=41'b00000011000010100001000100011011100000001;
1808:mir=41'b00000010000001100001000100010111100010010;
1809:mir=41'b10010100000000100101000111111000000101000;
40:mir=41'b10010100000000100101000111100000000000000;
41:mir=41'b10010100000000100101000111100000000000000;
42:mir=41'b10010100000000100101000111100000000000000;
43:mir=41'b10010100000000100101000111100000000000000;
44:mir=41'b10000100000001000000001010111011111111111;
1810:mir=41'b10010100000000100001000110000000000000000;
1811:mir=41'b00000011000010100001000100011011100010001;
1088:mir=41'b00000000000000000000000010111000000000010;
1116:mir=41'b00000000000000000000000010111000000000010;
2:mir=41'b10010100000000100001000101000000000000000;
3:mir=41'b10000100000000100001000111100000000000000;
4:mir=41'b10000100000000100001000111100000000000000;
5:mir=41'b10010100000000100101000111100000000000000;
6:mir=41'b10010100000000100101000111100000000000000;
7:mir=41'b10010100000000100101000111100000000000000;
8:mir=41'b10010101001010100101000100010100000001100;
9:mir=41'b10010101001010100101000100010100000001101;
10:mir=41'b10010101001010100101000100001000000001100;
11:mir=41'b00000000000000000000000010111011111111111;
12:mir=41'b10000001000010100000000100011000000000000;
13:mir=41'b10010101001010100101000100010100000010000;
14:mir=41'b00000000000000000000000010110000000001100;
15:mir=41'b00000000000000000000000010111011111111111;
16:mir=41'b00000000000000000000000010110100000010011;
17:mir=41'b00000000000000000000000010100100000001100;
18:mir=41'b00000000000000000000000010111011111111111;
19:mir=41'b00000000000000000000000010101100000001100;
20:mir=41'b00000000000000000000000010111011111111111;
2047:mir=41'b10000000000000100000000111011000000000000;

2046:mir=41'b11111111111111111111111111111111111111111;

default:mir=41'b10000001000000100101010010100000000000000;

endcase
end
	end
endmodule
