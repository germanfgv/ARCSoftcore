module decoder(
input[5:0] seleccion,
output reg [37:0] habilitador
);
initial habilitador=38'b0;

always@(seleccion)
begin
	habilitador[seleccion]=1'b1;
	case(seleccion)
		0:habilitador=38'b00000000000000000000000000000000000000;
		1:habilitador=38'b00000000000000000000000000000000000010;
		2:habilitador=38'b00000000000000000000000000000000000100;
		3:habilitador=38'b00000000000000000000000000000000001000;
		4:habilitador=38'b00000000000000000000000000000000010000;
		5:habilitador=38'b00000000000000000000000000000000100000;
		6:habilitador=38'b00000000000000000000000000000001000000;
		7:habilitador=38'b00000000000000000000000000000010000000;
		8:habilitador=38'b00000000000000000000000000000100000000;
		9:habilitador=38'b00000000000000000000000000001000000000;
		10:habilitador=38'b00000000000000000000000000010000000000;
		11:habilitador=38'b00000000000000000000000000100000000000;
		12:habilitador=38'b00000000000000000000000001000000000000;
		13:habilitador=38'b00000000000000000000000010000000000000;
		14:habilitador=38'b00000000000000000000000100000000000000;
		15:habilitador=38'b00000000000000000000001000000000000000;
		16:habilitador=38'b00000000000000000000010000000000000000;
		17:habilitador=38'b00000000000000000000100000000000000000;
		18:habilitador=38'b00000000000000000001000000000000000000;
		19:habilitador=38'b00000000000000000010000000000000000000;
		20:habilitador=38'b00000000000000000100000000000000000000;
		21:habilitador=38'b00000000000000001000000000000000000000;
		22:habilitador=38'b00000000000000010000000000000000000000;
		23:habilitador=38'b00000000000000100000000000000000000000;
		24:habilitador=38'b00000000000001000000000000000000000000;
		25:habilitador=38'b00000000000010000000000000000000000000;
		26:habilitador=38'b00000000000100000000000000000000000000;
		27:habilitador=38'b00000000001000000000000000000000000000;
		28:habilitador=38'b00000000010000000000000000000000000000;
		29:habilitador=38'b00000000100000000000000000000000000000;
		30:habilitador=38'b00000001000000000000000000000000000000;
		31:habilitador=38'b00000010000000000000000000000000000000;
		32:habilitador=38'b00000100000000000000000000000000000000;
		33:habilitador=38'b00001000000000000000000000000000000000;
		34:habilitador=38'b00010000000000000000000000000000000000;
		35:habilitador=38'b00100000000000000000000000000000000000;
		36:habilitador=38'b01000000000000000000000000000000000000;
		37:habilitador=38'b10000000000000000000000000000000000000;
		default:habilitador=38'b00000000000000000000000000000000000000;
	endcase
end
endmodule
